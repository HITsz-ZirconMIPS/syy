`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2021/07/02 22:37:43
// Design Name: 
// Module Name: data_ram
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


`include "defines.v"

module data_ram (
    input wire clk,
    input wire ce,
    input wire we,
    input wire[`DataAddrBus] raddr,
    input wire[`DataAddrBus] waddr,
    input wire[3:0] sel,
    input wire[`DataBus] data_i,

    output reg[`DataBus] data_o

);

wire[`DataAddrBus] addr = (ce)? raddr:(we)? waddr: `ZeroWord;

//定义四个字节数组(4个8位储存一个字)    DataMemNum 131071
reg [`ByteWidth] data_mem0[0:`DataMemNum-1] ;
reg [`ByteWidth] data_mem1[0:`DataMemNum-1] ;
reg [`ByteWidth] data_mem2[0:`DataMemNum-1] ;
reg [`ByteWidth] data_mem3[0:`DataMemNum-1] ;

//写操作 DataMemNumLog2为实际使用到的地址宽度，与 DataMemNum相对应
always @(posedge clk) begin
    if (ce == `ChipDisable) begin
        //data_o <= `ZeroWord;
    end else if (we == `WriteEnable) begin
        if (sel[3]==1'b1) begin
            data_mem3[addr[`DataMemNumLog2+1 : 2]] <= data_i[31:24];
        end
        if (sel[2]==1'b1) begin
            data_mem2[addr[`DataMemNumLog2+1 : 2]] <= data_i[24:16];
        end
        if (sel[1]==1'b1) begin
            data_mem1[addr[`DataMemNumLog2+1 : 2]] <= data_i[15:8];
        end
        if (sel[0]==1'b1) begin
            data_mem0[addr[`DataMemNumLog2+1 : 2]] <= data_i[7:0];
        end
        
    end
end

//读模块
always @(*) begin
    if (ce == `ChipDisable) begin
        data_o <= `ZeroWord;
    end else if (we == `WriteDisable) begin
        data_o <= {data_mem3[addr[`DataMemNumLog2+1 : 2]],
                    data_mem2[addr[`DataMemNumLog2+1 : 2]],
                    data_mem1[addr[`DataMemNumLog2+1 : 2]],
                    data_mem0[addr[`DataMemNumLog2+1 : 2]] };
    end else begin
        data_o <= `ZeroWord; 
    end
end

endmodule